----------------------------------------------------------------------------------
-- Company: CEM Solutions
-- Engineer: viru jawoor
-- 
-- Create Date:    17:30:26 05/20/2008 
-- Design Name:    RINGING TONE 
-- Module Name:    RAM- Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: SINE WAVE At 697Hz
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity iram_LUT is
    Port ( clk_5mhz : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           en : in  STD_LOGIC;
		   addr : in std_logic_vector(7 downto 0);
           ram_out : out  STD_LOGIC_vector(15 downto 0));
end iram_LUT;

architecture Behavioral of iram_LUT is

type ram is array  (0 to 204)of std_logic_vector (15 downto 0);
constant ram1 : ram :=(
-- "0010101010101101",
-- "0011101010111100",
-- "0010100100101001",
-- "0000011010001000",
-- "1110110010011101",
-- "1110100110111111",
-- "1111011100000001",
-- "0000000010110100",
-- "1111100101100000",
-- "1110011010010110",
-- "1101110001110100",
-- "1110101110001010",
-- "0001000010100010",
-- "0011010010110011",
-- "0011110111001100",
-- "0010001110001010",
-- "1111011001010010",
-- "1101001101000000",
-- "1100111001011011",
-- "1110010010001011",
-- "0000000001001111",
-- "0000110010001101",
-- "0000010110011100",
-- "1111101001101000",
-- "1111110101001010",
-- "0001001000011000",
-- "0010100100010110",
-- "0010101110101000",
-- "0001000000110001",
-- "1110010001001011",
-- "1100010000100111",
-- "1100010101111000",
-- "1110011011001110",
-- "0001000011101001",
-- "0010100011001011",
-- "0010001111100011",
-- "0000111000100100",
-- "1111110110111011",
-- "1111111101011101",
-- "0000101111110000",
-- "0001000000101100",
-- "1111111101000110",
-- "1110000001010110",
-- "1100101001111010",
-- "1101001001001101",
-- "1111100000000001",
-- "0010010100111101",
-- "0011110100011101",
-- "0011000110111100",
-- "0000111000001110",
-- "1110110001001010",
-- "1110000100001111",
-- "1110110001100001",
-- "1111110001100010",
-- "1111111010110111",
-- "1111000101010010",
-- "1110010000110110",
-- "1110101010101000",
-- "0000100010100111",
-- "0010110011011001",
-- "0011110011000111",
-- "0010100111100010",
-- "1111111000001101",
-- "1101010100001111",
-- "1100011111111000",
-- "1101101011011000",
-- "1111101101100010",
-- "0001000011110001",
-- "0001000001100100",
-- "0000001101101001",
-- "1111110110110001",
-- "0000100111101000",
-- "0001111100001110",
-- "0010011110100100",
-- "0001010011000000",
-- "1110110011001001",
-- "1100100011011011",
-- "1100001000110101",
-- "1101111010001000",
-- "0000101100100110",
-- "0010101100110001",
-- "0010110100111101",
-- "0001011100101011",
-- "1111111100000010",
-- "1111011101111101",
-- "0000000011001110",
-- "0000101000111110",
-- "0000001011000000",
-- "1110100111100000",
-- "1101001000011011",
-- "1101001000010101",
-- "1111000011100000",
-- "0001111000000001",
-- "0011110010000001",
-- "0011100010011001",
-- "0001011010000111",
-- "1110111011000000",
-- "1101101010100110",
-- "1110000110100001",
-- "1111010110101011",
-- "0000000101101101",
-- "1111101101110000",
-- "1110110111100111",
-- "1110110010100111",
-- "0000001000010101",
-- "0010001110111001",
-- "0011100011010011",
-- "0010111000001110",
-- "0000011000101000",
-- "1101100101111010",
-- "1100010001000100",
-- "1101000110110001",
-- "1111010001110100",
-- "0001001001111101",
-- "0001100111100010",
-- "0000110111000001",
-- "0000000011101100",
-- "0000001110100010",
-- "0001010001100001",
-- "0010000011101110",
-- "0001011011001111",
-- "1111010100010010",
-- "1100111111011000",
-- "1100000111011100",
-- "1101011101100110",
-- "0000001111010111",
-- "0010101010100101",
-- "0011010010110100",
-- "0010000011101000",
-- "0000001011110110",
-- "1111000111111010",
-- "1111010110111001",
-- "0000001000000010",
-- "0000001110000011",
-- "1111001010011000",
-- "1101101110001001",
-- "1101010011010010",
-- "1110101101100111",
-- "0001010110111101",
-- "0011100100000101",
-- "0011110100011001",
-- "0001111100010111",
-- "1111001110100101",
-- "1101011011111000",
-- "1101011110100010",
-- "1110110100100001",
-- "0000000101001101",
-- "0000010000011100",
-- "1111100011000111",
-- "1111000101111010",
-- "1111110110011010",
-- "0001101000101100",
-- "0011001000111111",
-- "0010111110001111",
-- "0000110111000011",
-- "1101111111111100",
-- "1100001110000010",
-- "1100100111101100",
-- "1110110000111011",
-- "0001000100101101",
-- "0010000101011100",
-- "0001100010011100",
-- "0000011010111011",
-- "1111111111010001",
-- "0000100111110010",
-- "0001100000000011",
-- "0001011000001011",
-- "1111110001001001",
-- "1101100001110001",
-- "1100010001111111",
-- "1101001000101011",
-- "1111101111001000",
-- "0010011101010111",
-- "0011100110101110",
-- "0010101001111010",
-- "0000100100101010",
-- "1110111100111000",
-- "1110101110010011",
-- "1111100000011010",
-- "0000000101101100",
-- "1111100110110010",
-- "1110010111111010",
-- "1101101001100010",
-- "1110100000111001",
-- "0000110101001110",
-- "0011001100000110",
-- "0011111011001110",
-- "0010011011011111",
-- "1111101001100100",
-- "1101011000111001",
-- "1100111100110110",
-- "1110001110000100",
-- "1111111001100111",
-- "0000101010101001",
-- "0000001111111100",
-- "1111100011010001",
-- "1111101110110010",
-- "0001000100010010",
-- "0010100110010010",
-- "0010111000100010",
-- "0001010000001000",
-- "1110011111011100",
-- "1100010110110110",
-- "1100010001000010",
-- "1110001110001010");   -------Key1  P2P2b4V 

-- "0101100011001110",
-- "0111000000101110",
-- "0011111101101111",
-- "1111110001110000",
-- "1110001000011001",
-- "1111011110110000",
-- "0000111100100010",
-- "1111101001100110",
-- "1100000001000010",
-- "1001100110011100",
-- "1011100011000111",
-- "0001001110101000",
-- "0110011110100101",
-- "0111010101010000",
-- "0011100111110010",
-- "1110111100010100",
-- "1101000101010010",
-- "1110011111001101",
-- "0000001110100011",
-- "1111011000011100",
-- "1100010100001000",
-- "1010011100110000",
-- "1100101110111101",
-- "0010010111011001",
-- "0111001010011100",
-- "0111010101001111",
-- "0010111110011000",
-- "1101111010001010",
-- "1011111111110110",
-- "1101101000010011",
-- "1111110001101001",
-- "1111011011111001",
-- "1100111001011100",
-- "1011011101100110",
-- "1101111010011011",
-- "0011010100111010",
-- "0111100011011100",
-- "0111000000011010",
-- "0010000100010110",
-- "1100110000011101",
-- "1010111110000001",
-- "1100111110111111",
-- "1111101000011000",
-- "1111110011011011",
-- "1101101101011110",
-- "1100100011011110",
-- "1110111111101011",
-- "0100000010101100",
-- "0111100111110011",
-- "0110011000001010",
-- "0000111101111000",
-- "1011100100111100",
-- "1010000101011010",
-- "1100100111001011",
-- "1111110011110000",
-- "0000011100110010",
-- "1110101011011100",
-- "1101101000011111",
-- "1111111001011010",
-- "0100011101100010",
-- "0111010111011001",
-- "0101011111011101",
-- "1111110000001101",
-- "1010011101100010",
-- "1001011010111011",
-- "1100100011010010",
-- "0000010011000011",
-- "0001010100010111",
-- "1111101101110100",
-- "1110100110110100",
-- "0000100011001101",
-- "0100100011110011",
-- "0110110011101111",
-- "0100011010100110",
-- "1110100001000110",
-- "1001011111110100",
-- "1001000010010101",
-- "1100110100001001",
-- "0001000011111010",
-- "0010010101010010",
-- "0000101110101101",
-- "1111011001001110",
-- "0000111010000010",
-- "0100010101011101",
-- "0101111111111011",
-- "0011001110110110",
-- "1101010110011101",
-- "1000110000101000",
-- "1000111101111101",
-- "1101011000111010",
-- "0010000010100101",
-- "0011011001111111",
-- "0001101000010100",
-- "1111111011011011",
-- "0000111100010101",
-- "0011110100001110",
-- "0101000000010111",
-- "0010000010000010",
-- "1100010101110111",
-- "1000010011100111",
-- "1001001110011101",
-- "1110001111000110",
-- "0011001010001000",
-- "0100011100100010",
-- "0010010101011111",
-- "0000001010011101",
-- "0000101010010001",
-- "0011000011010001",
-- "0011111010010110",
-- "0000111010000010",
-- "1011100100000001",
-- "1000001010111100",
-- "1001110010111000",
-- "1111010010110101",
-- "0100010100111011",
-- "0101010111001101",
-- "0010110010000000",
-- "0000000100111101",
-- "0000000101101010",
-- "0010000111000110",
-- "0010110011110000",
-- "1111111100010111",
-- "1011000100011110",
-- "1000010111001100",
-- "1010101000100101",
-- "0000011111000111",
-- "0101011101000010",
-- "0110000100110111",
-- "0010111011000101",
-- "1111101011001110",
-- "1111010001110101",
-- "0001000101000101",
-- "0001110010011011",
-- "1111001101101010",
-- "1010111001010011",
-- "1000110111001110",
-- "1011101011100101",
-- "0001101110001111",
-- "0110011100110001",
-- "0110100001011100",
-- "0010101111011101",
-- "1110111111001101",
-- "1110010011010110",
-- "0000000011000101",
-- "0000111011110100",
-- "1110110001010110",
-- "1011000010111000",
-- "1001101000010010",
-- "1100110110110100",
-- "0010111010010010",
-- "0111001111000010",
-- "0110101010010000",
-- "0010001111100110",
-- "1110000100010110",
-- "1101001111101011",
-- "1111000110111101",
-- "0000010100011110",
-- "1110101001010110",
-- "1011011111111101",
-- "1010100110010011",
-- "1110000100100011",
-- "0011111101100110",
-- "0111101111111010",
-- "0110011110001100",
-- "0001011101100110",
-- "1100111111010101",
-- "1100001100101011",
-- "1110010110000110",
-- "1111111111101101",
-- "1110110101111010",
-- "1100001101101100",
-- "1011101100001000",
-- "1111001110110111",
-- "0100110011001011",
-- "0111111100110011",
-- "0101111101110111",
-- "0000011101000000",
-- "1011110101101001",
-- "1011010000001011",
-- "1101110100111011",
-- "1111111111010010",
-- "1111010101101000",
-- "1101000111110110",
-- "1100110011111111",
-- "0000010000001000",
-- "0101010111001011",
-- "0111110100110000",
-- "0101001011011101",
-- "1111010010100101",
-- "1010101101001101",
-- "1010011111100000",
-- "1101100110101001",
-- "0000010011010100",
-- "0000000101100010",
-- "1110001001010000",
-- "1101111000000000",
-- "0001000011011100",
-- "0101100111001001",
-- "0111011000100000",
-- "0100001010101100",
-- "1110000011111010",
-- "1001101011110011",
-- "1001111111000001",
-- "1101101100110111",
-- "0000111010010000"); --key2

-- "0101101111111101",
-- "0110011110111111",
-- "0010101010010101",
-- "1111010001001100",
-- "1111101101110110",
-- "0001111011111010",
-- "0001010011111101",
-- "1100110010111100",
-- "1000101100010101",
-- "1001110100001011",
-- "1111101111001010",
-- "0101000010001101",
-- "0101010011110011",
-- "0001111001011011",
-- "1111110001101110",
-- "0001010101001101",
-- "0011100010001000",
-- "0001111010111011",
-- "1100011111010001",
-- "1000010000110100",
-- "1001101100110011",
-- "1111100000111110",
-- "0100000110001011",
-- "0011110110000100",
-- "0000111100010010",
-- "0000001011011111",
-- "0010110100100011",
-- "0100111110111100",
-- "0010100000100001",
-- "1100011010100000",
-- "1000001111101011",
-- "1001111011011001",
-- "1111010111110110",
-- "0011000000000111",
-- "0010001010111001",
-- "1111110101110111",
-- "0000011101000010",
-- "0100000110111000",
-- "0110001100111000",
-- "0011000001011001",
-- "1100100011011110",
-- "1000101000100110",
-- "1010100000001001",
-- "1111010101101111",
-- "0001110100101011",
-- "0000011000001000",
-- "1110101001111011",
-- "0000100101110011",
-- "0101001000000101",
-- "0111000111010001",
-- "0011011010010001",
-- "1100111000001000",
-- "1001011001110001",
-- "1011011001111010",
-- "1111011011111110",
-- "0000101000100110",
-- "1110100100000100",
-- "1101011100110101",
-- "0000100110000011",
-- "0101110101001111",
-- "0111101010011100",
-- "0011101000010000",
-- "1101010101110000",
-- "1010100000000011",
-- "1100100110001101",
-- "1111101011000111",
-- "1111100000011000",
-- "1100110101000111",
-- "1100010011010010",
-- "0000011110110101",
-- "0110001100101010",
-- "0111110100000011",
-- "0011101001000000",
-- "1101111001001111",
-- "1011110111000111",
-- "1110000001010110",
-- "0000000010110101",
-- "1110100000000000",
-- "1011010001010101",
-- "1011010010000011",
-- "0000010001111011",
-- "0110001110000001",
-- "0111100011001010",
-- "0011011010111111",
-- "1110011111001111",
-- "1101011001110011",
-- "1111100110101000",
-- "0000100001111111",
-- "1101101010101110",
-- "1001111110001001",
-- "1010011101100111",
-- "0000000001100110",
-- "0101111010010011",
-- "0110111000011010",
-- "0010111101101011",
-- "1111000100100000",
-- "1111000010010110",
-- "0001010000101000",
-- "0001000110101001",
-- "1101000010110101",
-- "1000111111111111",
-- "1001111001110111",
-- "1111110000011101",
-- "0101010011101101",
-- "0101110101110111",
-- "0010010001100010",
-- "1111100110000111",
-- "0000101010110111",
-- "0010111001011101",
-- "0001101110001011",
-- "1100101001101001",
-- "1000011010000101",
-- "1001101001110110",
-- "1111100001001011",
-- "0100011101011011",
-- "0100011111000010",
-- "0001011000001011",
-- "0000000001101011",
-- "0010001101100100",
-- "0100011011001010",
-- "0010010101100000",
-- "1100011111010111",
-- "1000001110001100",
-- "1001101111100010",
-- "1111010110010001",
-- "0011011011100000",
-- "0010111000100110",
-- "0000010100001011",
-- "0000010101100000",
-- "0011100101001100",
-- "0101110000000100",
-- "0010111001010001",
-- "1100100011001010",
-- "1000011100100111",
-- "1010001011100110",
-- "1111010001111001",
-- "0010010010011100",
-- "0001001000001001",
-- "1111001001000011",
-- "0000100000110000",
-- "0100101101010010",
-- "0110110011000111",
-- "0011010110000110",
-- "1100110011010110",
-- "1001000100001000",
-- "1010111101011011",
-- "1111010101100101",
-- "0001000110111011",
-- "1111010011110110",
-- "1101111011000000",
-- "0000100011011000",
-- "0101100010011110",
-- "0111100000001101",
-- "0011101000111010",
-- "1101001101011011",
-- "1010000010000101",
-- "1100000011000010",
-- "1111100010001011",
-- "1111111101100011",
-- "1101100010000110",
-- "1100101110101011",
-- "0000011110001101",
-- "0110000010100010",
-- "0111110100011101",
-- "0011101111000110",
-- "1101101110011010",
-- "1011010010100111",
-- "1101011001001010",
-- "1111110111101001",
-- "1110111010100000",
-- "1011111001001010",
-- "1011101000110111",
-- "0000010010110000",
-- "0110001100101011",
-- "0111101110010110",
-- "0011100110110100",
-- "1110010011000100",
-- "1100110000110111",
-- "1110111011011101",
-- "0000010101001001",
-- "1110000001010100",
-- "1010011110101110",
-- "1010101110001111",
-- "0000000011001010",
-- "0110000001010101",
-- "0111001101111000",
-- "0011001111001000",
-- "1110111000000101",
-- "1110010111010010",
-- "0000100100101111",
-- "0000111000111101",
-- "1101010100100111",
-- "1001010111101010",
-- "1010000010111111",
-- "1111110001111100",
-- "0101100010010001",
-- "0110010100100110",
-- "0010101000001001",
-- "1111011010011011",
-- "0000000000000000",
-- "0010001111001111",
-- "0001100000101011",
-- "1100110110000100",
-- "1000100111101011",
-- "1001101010100010");  -------Key3



-- "0101100001101110",
-- "0111100001110011",
-- "0101000010011000",
-- "0000001101000010",
-- "1100011110010000",
-- "1011111010101010",
-- "1101110111111000",
-- "1111111001100101",
-- "0000000110011100",
-- "1110110010001010",
-- "1110000010001101",
-- "1111100111110110",
-- "0011000111100100",
-- "0101111011101001",
-- "0101010111001011",
-- "0000111110011110",
-- "1011010010111011",
-- "1000000110000000",
-- "1001100101100111",
-- "1110101111110110",
-- "0100000101001011",
-- "0110010000100101",
-- "0100100000000011",
-- "0000110110110000",
-- "1110010010001110",
-- "1110001101111001",
-- "1111100111000001",
-- "0000001101011010",
-- "1110110100101100",
-- "1100100011110111",
-- "1011111011000011",
-- "1110011111110011",
-- "0011010000010100",
-- "0111000000111001",
-- "0110110100001100",
-- "0010010101010110",
-- "1100010100100001",
-- "1000101010010011",
-- "1001100001101111",
-- "1101111000010100",
-- "0010011100101010",
-- "0100010101001111",
-- "0011000110100101",
-- "0000110000001111",
-- "1111101100001101",
-- "0000100100001101",
-- "0001110100001000",
-- "0001010000101011",
-- "1110010101011110",
-- "1010111010111000",
-- "1001111110010001",
-- "1101000001010001",
-- "0010100111100100",
-- "0111001010111111",
-- "0111100011010010",
-- "0011011110001010",
-- "1101101101110111",
-- "1010000010010110",
-- "1010011000110101",
-- "1101101100100000",
-- "0001000001110100",
-- "0010000110111111",
-- "0001000010010110",
-- "1111110110010010",
-- "0000011010010111",
-- "0010100011011111",
-- "0100000110011110",
-- "0010110101000010",
-- "1110101001111011",
-- "1010000111001110",
-- "1000100100101011",
-- "1011100100111100",
-- "0001011101010111",
-- "0110011011111110",
-- "0111010111111100",
-- "0100000010001111",
-- "1111000101101110",
-- "1011111011000111",
-- "1100000100110001",
-- "1110010101101101",
-- "0000001010010101",
-- "0000000000010100",
-- "1110101001000001",
-- "1110010001101110",
-- "0000010101010100",
-- "0011110110111101",
-- "0110000011100001",
-- "0100100011111100",
-- "1111100111011010",
-- "1010001101101000",
-- "1000000000011011",
-- "1010100011110110",
-- "0000001000111101",
-- "0101000001011100",
-- "0110010001011101",
-- "0011110010101000",
-- "0000000011111011",
-- "1101111011011110",
-- "1110010100011111",
-- "1111110001001111",
-- "0000000011001111",
-- "1110011001010110",
-- "1100010101000000",
-- "1100010101100100",
-- "1111100001110101",
-- "0100010011100101",
-- "0111010100101101",
-- "0110000011100000",
-- "0000111001111001",
-- "1011000110101001",
-- "1000011000111111",
-- "1010010001110000",
-- "1111000011101011",
-- "0011010001100110",
-- "0100011011001010",
-- "0010101011100110",
-- "0000010110101000",
-- "1111101001101000",
-- "0000101111011101",
-- "0001110000111011",
-- "0000101101111011",
-- "1101100010101000",
-- "1010011111110101",
-- "1010011010111001",
-- "1110001111100010",
-- "0011111010001111",
-- "0111101100001110",
-- "0110111100010001",
-- "0010001000011011",
-- "1100100000011010",
-- "1001101001101000",
-- "1010111000110001",
-- "1110100011001001",
-- "0001100110010011",
-- "0010001001111110",
-- "0000110101011111",
-- "1111110110010011",
-- "0000110000101001",
-- "0010111010111101",
-- "0011111110000001",
-- "0010000000000001",
-- "1101100001101100",
-- "1001011100101100",
-- "1000111011011110",
-- "1100110101100111",
-- "0010110111011111",
-- "0111000111111001",
-- "0110111110010011",
-- "0010111010110001",
-- "1110000010100111",
-- "1011100010011001",
-- "1100010111000000",
-- "1110110100100100",
-- "0000010111011000",
-- "1111111000000010",
-- "1110100011001010",
-- "1110100111011111",
-- "0001000101000100",
-- "0100011111101111",
-- "0101111110000111",
-- "0011100101011111",
-- "1110001111111100",
-- "1001010100011100",
-- "1000001100001010",
-- "1011101101011111",
-- "0001100000101010",
-- "0101110001101100",
-- "0110000100110000",
-- "0010111110110100",
-- "1111010011111010",
-- "1101101011100010",
-- "1110011110110101",
-- "1111111001101000",
-- "1111110101100010",
-- "1101111111000001",
-- "1100001101111010",
-- "1100111001110100",
-- "0000100111001101",
-- "0101001110111100",
-- "0111011000110010",
-- "0101000101001100",
-- "1111011100010001",
-- "1010000011101101",
-- "1000011000010010",
-- "1011001101001111",
-- "0000001111000011",
-- "0011111101011101",
-- "0100010111000001",
-- "0010001100100111",
-- "1111111111100010",
-- "1111101010101001",
-- "0000111001110010",
-- "0001101000000100",
-- "0000000110100101",
-- "1100110010101111",
-- "1010010000001001",
-- "1011000100101001",
-- "1111100011000100",
-- "0101000101001101",
-- "0111111100110110",
-- "0110000110010101",
-- "0000101110111000",
-- "1011011011110010",
-- "1001011111010000",
-- "1011100010101100");---key4

-- "0101101111100001",
-- "0111001100101001",
-- "0011110110110110",
-- "1111001010100010",
-- "1101000001101111",
-- "1110001011011011",
-- "1111111100011000",
-- "1111011101100011",
-- "1100111100011111",
-- "1011100011111010",
-- "1110000001101011",
-- "0011011010001011",
-- "0111100001000110",
-- "0110101011010011",
-- "0001010000100100",
-- "1011011110011110",
-- "1001100101101001",
-- "1100001011001100",
-- "0000000001010101",
-- "0001100011111011",
-- "0000010110110101",
-- "1111001000111011",
-- "0000100010000111",
-- "0011111010111001",
-- "0101110010010101",
-- "0011010010011001",
-- "1101011100101100",
-- "1000101010010100",
-- "1000110011000010",
-- "1101101001110100",
-- "0011001011011101",
-- "0101001111111110",
-- "0011010011010101",
-- "0000010111001101",
-- "1111101000010000",
-- "0001001011001000",
-- "0010000110110110",
-- "1111111100110111",
-- "1011101011001100",
-- "1001001001010000",
-- "1011011001010001",
-- "0001011010000011",
-- "0110101100010010",
-- "0111001111110110",
-- "0011000111010001",
-- "1110000111101001",
-- "1100001001111001",
-- "1101101010011101",
-- "1111101111011001",
-- "1111100010100110",
-- "1101011001110110",
-- "1100011101101111",
-- "1111001001111100",
-- "0100001111000110",
-- "0111100001010101",
-- "0101110000011000",
-- "1111110111100110",
-- "1010010101100101",
-- "1001001100111111",
-- "1100100011001111",
-- "0000110010111110",
-- "0010010111010110",
-- "0001000010001001",
-- "1111101011010101",
-- "0000110101100001",
-- "0011110000000000",
-- "0100111110011100",
-- "0010000001111000",
-- "1100010100100111",
-- "1000010010110001",
-- "1001011010010110",
-- "1110111001011101",
-- "0100011000101001",
-- "0101111001011100",
-- "0011010011000010",
-- "1111111011110000",
-- "1111000001001101",
-- "0000011101100101",
-- "0001010100011101",
-- "1111010001110010",
-- "1011011111100001",
-- "1001101111101000",
-- "1100101001101101",
-- "0010101111001000",
-- "0111011001010110",
-- "0110111111011000",
-- "0010001000000011",
-- "1100111110100100",
-- "1011010110010110",
-- "1101010101101100",
-- "1111110010010101",
-- "1111110110110100",
-- "1110000001010000",
-- "1101011000110100",
-- "0000001001000001",
-- "0100110010101000",
-- "0111001110010010",
-- "0100101000010100",
-- "1110011101010100",
-- "1001010111100001",
-- "1001000110010010",
-- "1101001100111101",
-- "0001101111111011",
-- "0011001100111000",
-- "0001100110101001",
-- "0000000000001111",
-- "0000111000011000",
-- "0011010110010100",
-- "0100000010111111",
-- "0000110100110111",
-- "1011011010111000",
-- "1000001111001010",
-- "1010010010111001",
-- "0000010000100010",
-- "0101100001000001",
-- "0110010100110000",
-- "0011000001010000",
-- "1111010001100001",
-- "1110010010000101",
-- "1111110000100100",
-- "0000101011001101",
-- "1110110110011100",
-- "1011100101100100",
-- "1010100011001100",
-- "1101111100111011",
-- "0011111010100111",
-- "0111110100000101",
-- "0110011011100001",
-- "0000111100010000",
-- "1011110011111101",
-- "1010101011101001",
-- "1101010000000011",
-- "0000000101100001",
-- "0000010111111000",
-- "1110101110100010",
-- "1110010000011100",
-- "0000111011010101",
-- "0101000011101001",
-- "0110101001110100",
-- "0011010111010011",
-- "1101000110101011",
-- "1000101000001010",
-- "1001010010111001",
-- "1110000110110011",
-- "0010110100010110",
-- "0011111111110100",
-- "0010000000010110",
-- "0000000101101100",
-- "0000101011011000",
-- "0010110001000101",
-- "0011000100101001",
-- "1111101111111001",
-- "1010110010001101",
-- "1000011111010001",
-- "1011011001100111",
-- "0001101010010000",
-- "0110011111111001",
-- "0110011111000001",
-- "0010011101110111",
-- "1110011011000000",
-- "1101011111001010",
-- "1111001000101010",
-- "0000001110011111",
-- "1110101011110100",
-- "1011111011100001",
-- "1011011111111000",
-- "1111001110000001",
-- "0100111000100100",
-- "0111111010111111",
-- "0101100101110110",
-- "1111100111111000",
-- "1010101100101100",
-- "1010001101110010",
-- "1101011011010001",
-- "0000100111111111",
-- "0001000010011101",
-- "1111011101000100",
-- "1111000000010000",
-- "0001011110010010",
-- "0101000010010110",
-- "0101110110111001",
-- "0010000010000101",
-- "1011111000011111",
-- "1000001010011111",
-- "1001110010111011",
-- "1111001110000001",
-- "0011111011110001",
-- "0100101011100010",
-- "0010001100000011",
-- "1111111010111101",
-- "0000010000011101",
-- "0010000100010010",
-- "0010001000001011",
-- "1110110110110100",
-- "1010011100000111",
-- "1001000001100111",
-- "1100101010100001",
-- "0011000001101001",
-- "0111010001001001",
-- "0110010110011110",
-- "0001101001111111",
-- "1101011011110010",
-- "1100101101000111",
-- "1110101010000011",
-- "0000000000101001");--key5




"0101111100010000",
"0110101010111010",
"0010100011011100",
"1110101001111110",
"1110100111001100",
"0000101000100101",
"0000010011110011",
"1100100110111001",
"1001100111110001",
"1011110001101001",
"0010001101101110",
"0111001101101111",
"0110010110010011",
"0001001111011111",
"1101011010100000",
"1101110111011000",
"0000000010011111",
"1111100110111010",
"1100010010000011",
"1010011100010100",
"1101101111100000",
"0100001101001001",
"0111111001010101",
"0101011001100100",
"1111100100001011",
"1100001000101001",
"1101010010110111",
"1111101111000101",
"1111010011101100",
"1100011100000010",
"1011101001011111",
"1111101111011101",
"0101110001101110",
"0111111001101101",
"0011111000101110",
"1101101100000110",
"1011000000011100",
"1101000011010101",
"1111110011101111",
"1111011010001100",
"1100111110101110",
"1101000011101001",
"0001100100000011",
"0110110010001011",
"0111001110011110",
"0001111100010010",
"1011110100001001",
"1010001101100101",
"1101001111101010",
"0000010001101110",
"1111110110001111",
"1101110000111011",
"1110011110010011",
"0011000001110101",
"0111001001100011",
"0101111100001100",
"1111110000001111",
"1010001001111011",
"1001111001101001",
"1101111010111100",
"0001000110000010",
"0000100000001010",
"1110100111101101",
"1111101101110110",
"0100000000110100",
"0110110111110101",
"0100001011110001",
"1101100010101000",
"1000111010000101",
"1010001010110010",
"1111000011110011",
"0010001001101110",
"0001001101111010",
"1111011000000110",
"0000101001000100",
"0100011101010010",
"0110000001101100",
"0010001001011100",
"1011100001110111",
"1000001110100011",
"1011000010101111",
"0000100100011011",
"0011010010110101",
"0001110100101010",
"1111111000101010",
"0001001010010101",
"0100011000001110",
"0100101111111011",
"0000000011000111",
"1001111010111011",
"1000001101010111",
"1100011110011011",
"0010010011001111",
"0100010101110011",
"0010001010010110",
"0000000010111010",
"0001010000010010",
"0011110110111010",
"0011001110000110",
"1110000110110000",
"1000110111110100",
"1000110111101110",
"1110010110010000",
"0100000100000010",
"0101000111000010",
"0010000111010100",
"1111110100001101",
"0000111101111011",
"0011000010000110",
"0001101001000000",
"1100100000100001",
"1000011110010010",
"1010001001111000",
"0000011110111000",
"0101101001100001",
"0101011100100101",
"0001100111011011",
"1111001110001110",
"0000011001111110",
"0010000100101000",
"0000001100111110",
"1011011001011011",
"1000101111010010",
"1011111011100010",
"0010101010101000",
"0110110111000001",
"0101001111101001",
"0000101010110101",
"1110010110101100",
"1111101101111011",
"0001001001111000",
"1111000100001111",
"1010110110010000",
"1001100110110101",
"1110000000110101",
"0100101011000111",
"0111100010001011",
"0100011101100100",
"1111010110000111",
"1101010110100110",
"1111000100100000",
"0000011100000100",
"1110010101101001",
"1010110111000011",
"1010111100101010",
"0000001011111001",
"0110010011000011",
"0111100100010101",
"0011001000011001",
"1101110001110011",
"1100011000111111",
"1110101000000110",
"0000000010110100",
"1110000011110100",
"1011010111010111",
"1100100101011000",
"0010001110011100",
"0111010111110110",
"0110111011011101",
"0001010110110100",
"1100001001010010",
"1011101001010001",
"1110100001001000",
"0000000010000101",
"1110001101000001",
"1100001110111110",
"1110010011111101",
"0011111011101000",
"0111110010111100",
"0101101010011101",
"1111010011010110",
"1010101001011100",
"1011010001101010",
"1110110100110001",
"0000011001100010",
"1110101011011010",
"1101010011001000",
"1111111011011110",
"0101001001100101",
"0111100010100011",
"0011111000111011",
"1101001011001011",
"1001011110111000",
"1011011001101010",
"1111100100001000",
"0001000100101111",
"1111010110001001",
"1110011000001001",
"0001010000101111",
"0101110010011111",
"0110101001111001",
"0001110010010000",
"1011001100100001",
"1000110100010001",
"1100000100110011",
"0000101011110111",
"0001111011101010",
"0000000010101001",
"1111010011000100",
"0010001011110010",
"0101110101010100",
"0101010000101010",
"1111100100001011",
"1001100100110111",
"1000110000111010");--key6

-- "0101101110111110",
-- "0111101011011100",
-- "0100110001111010",
-- "1111010110100001",
-- "1011001100010000",
-- "1010101110001110",
-- "1101011011001010",
-- "0000101010010110",
-- "0010000011001000",
-- "0001010011100110",
-- "0000000111010100",
-- "0000010000001010",
-- "0001110001011110",
-- "0010111000101011",
-- "0001101011010111",
-- "1110001000110000",
-- "1010100110100011",
-- "1010000100111011",
-- "1101101100100100",
-- "0011011110101100",
-- "0111100010001011",
-- "0110111001110011",
-- "0001110110100010",
-- "1011110000011111",
-- "1000101001101101",
-- "1010010011101111",
-- "1111000111011010",
-- "0011100001011000",
-- "0100110011010001",
-- "0010111010111111",
-- "0000000111110110",
-- "1110110000010110",
-- "1111010100000001",
-- "0000010011000010",
-- "1111111010110001",
-- "1110000000010101",
-- "1100010111001001",
-- "1101001010110001",
-- "0000110100000010",
-- "0101000110111011",
-- "0110101111111001",
-- "0011111100111010",
-- "1110000111111111",
-- "1001000101110010",
-- "1000010101111011",
-- "1100011011110011",
-- "0010100011000010",
-- "0110100101100100",
-- "0110001010101111",
-- "0010001011011111",
-- "1101110011111100",
-- "1011111100101011",
-- "1101000101101100",
-- "1111011000110011",
-- "0000100101000111",
-- "0000000001100100",
-- "1111000101011111",
-- "1111100110101110",
-- "0001111001111100",
-- "0100001100100010",
-- "0100000000101011",
-- "0000100000100011",
-- "1011100110110001",
-- "1000110011110101",
-- "1010100010110001",
-- "0000000101001010",
-- "0101110110000000",
-- "0111111100001001",
-- "0101000000111110",
-- "1111001101110111",
-- "1010100001100100",
-- "1001110011001011",
-- "1100110110010110",
-- "0000111011110000",
-- "0011001000110010",
-- "0010100101110110",
-- "0000110001111110",
-- "1111110110111011",
-- "0000100100011110",
-- "0001101001000110",
-- "0001001000111001",
-- "1110100001110101",
-- "1011100010100001",
-- "1010111010001101",
-- "1101111111110000",
-- "0011010010000011",
-- "0111001011111000",
-- "0110101100010111",
-- "0001110001011001",
-- "1011100101100110",
-- "1000010001001000",
-- "1001111001101011",
-- "1111000101100110",
-- "0100000111110110",
-- "0101110100101101",
-- "0011101111101111",
-- "0000001000100100",
-- "1101110100110101",
-- "1101111101011000",
-- "1111010111001010",
-- "1111111111010010",
-- "1111000000100001",
-- "1101101000010010",
-- "1101111011001001",
-- "0000101100101010",
-- "0100010111001111",
-- "0101111100111001",
-- "0011100011011000",
-- "1110001010100000",
-- "1001010010100101",
-- "1000011100100001",
-- "1100011101010100",
-- "0010101110010100",
-- "0111000011111001",
-- "0110101111111100",
-- "0010011010100000",
-- "1101010110001010",
-- "1010111001001110",
-- "1100000011000111",
-- "1111000100100100",
-- "0001010001111101",
-- "0001010111000101",
-- "0000001110110111",
-- "1111110110110110",
-- "0001001010000111",
-- "0010111111001000",
-- "0011000110110110",
-- "0000010111110101",
-- "1100001000100001",
-- "1001100000110001",
-- "1010111110011101",
-- "0000001001110110",
-- "0101110001111011",
-- "0111111101110001",
-- "0101000110001011",
-- "1111000110000001",
-- "1010000000101110",
-- "1001000100000010",
-- "1100011000100101",
-- "0001001100110011",
-- "0100001001010101",
-- "0011110010110010",
-- "0001011001100111",
-- "1111011100010000",
-- "1111010101100110",
-- "0000010110111111",
-- "0000100101110010",
-- "1110111111001010",
-- "1100100111011101",
-- "1011111000100110",
-- "1110010101101110",
-- "0010111110011100",
-- "0110100111110010",
-- "0110010010011100",
-- "0001101001000100",
-- "1011100010111110",
-- "1000000111001001",
-- "1001101011100001",
-- "1111000110010100",
-- "0100100111010011",
-- "0110101011001101",
-- "0100011100011101",
-- "0000000111011110",
-- "1100111100010001",
-- "1100101010101000",
-- "1110011101110010",
-- "0000000101100110",
-- "0000000011101111",
-- "1110111101101111",
-- "1110101110001010",
-- "0000100010011110",
-- "0011011110100010",
-- "0100111110110110",
-- "0011000011111101",
-- "1110010001001101",
-- "1001101100010101",
-- "1000110001011000",
-- "1100100101100010",
-- "0010110100101010",
-- "0111010101000001",
-- "0111001000000110",
-- "0010100100000100",
-- "1100111100010111",
-- "1001111111000001",
-- "1011001000101111",
-- "1110110011101001",
-- "0001111101110101",
-- "0010101010011010",
-- "0001010110110011",
-- "0000000101011110",
-- "0000010110101100",
-- "0001101011110111",
-- "0010001000000111",
-- "0000001111110100",
-- "1100110010100000",
-- "1010011010000001",
-- "1011100011000101",
-- "0000001101101001",
-- "0101100010101001",
-- "0111110000010100",
-- "0101000001101000",
-- "1110111111100000",
-- "1001101010110101",
-- "1000100010001100",
-- "1100000010100011");--KEY7 2v


-- "0101111100110010",
-- "0111010110010010",
-- "0011100110011000",
-- "1110010100000001",
-- "1011101111101111",
-- "1100111111000000",
-- "1111011111101010",
-- "0000001110010101",
-- "1110111001001011",
-- "1110000101010101",
-- "0000000110110011",
-- "0100000010011111",
-- "0110001011000000",
-- "0011101000010101",
-- "1101100100110000",
-- "1000101000110000",
-- "1000111001010001",
-- "1110001010000111",
-- "0100001000010010",
-- "0110010010110001",
-- "0011110011110101",
-- "1111110010001010",
-- "1101111000100110",
-- "1110110100101001",
-- "0000001001110101",
-- "1111011000001111",
-- "1100111101000101",
-- "1011111110010010",
-- "1110110001100111",
-- "0100000000111100",
-- "0111011000010000",
-- "0101100000100001",
-- "1111010111000010",
-- "1001101001010110",
-- "1000101110110101",
-- "1100110110001000",
-- "0010001001011101",
-- "0100011101010101",
-- "0010111101011111",
-- "0000010111110111",
-- "1111101100100001",
-- "0001000001101110",
-- "0001101101101100",
-- "1111100101011010",
-- "1011110000111111",
-- "1001111111001111",
-- "1100111000110011",
-- "0010111111010110",
-- "0111100100101010",
-- "0110110011001101",
-- "0001001111100001",
-- "1011011001001010",
-- "1001101000000100",
-- "1100011100111001",
-- "0000100011001010",
-- "0010010011110010",
-- "0001001111001111",
-- "1111111001111101",
-- "0000101110000111",
-- "0011000011010001",
-- "0011110001110101",
-- "0000110000111010",
-- "1011100110100100",
-- "1000101000111000",
-- "1010111101111100",
-- "0001010001101010",
-- "0110101101111111",
-- "0111001000111110",
-- "0010101011101010",
-- "1101011001011010",
-- "1011010111001111",
-- "1101000111101100",
-- "1111110001101001",
-- "0000011001001110",
-- "1111000011111000",
-- "1110011111011000",
-- "0000101101011100",
-- "0100011001011001",
-- "0101110100001001",
-- "0010100101001011",
-- "1100011110000100",
-- "1000010001001001",
-- "1001100011001101",
-- "1111010111100111",
-- "0101000011110010",
-- "0110011010011110",
-- "0011010000011001",
-- "1111000111000000",
-- "1101100000010110",
-- "1110101101101010",
-- "0000000011000010",
-- "1111001100101001",
-- "1100111101111001",
-- "1100011111001110",
-- "1111101100010001",
-- "0100101111101110",
-- "0111010010111011",
-- "0100100001101011",
-- "1110000110001101",
-- "1000111101011011",
-- "1001000010010101",
-- "1101110100001001",
-- "0011000011001101",
-- "0100110010011101",
-- "0010110001011110",
-- "0000000011111010",
-- "1111100000100011",
-- "0000110110001101",
-- "0001010011100111",
-- "1111000000110010",
-- "1011011110011011",
-- "1010011010101110",
-- "1101111101100011",
-- "0100000010110100",
-- "0111110101110011",
-- "0110000011101010",
-- "0000000000110010",
-- "1010100001000111",
-- "1001100101101111",
-- "1101000100001101",
-- "0001001111001111",
-- "0010101010111001",
-- "0001010100100110",
-- "1111111111001001",
-- "0000110111100000",
-- "0010111111100001",
-- "0011001110101110",
-- "1111110111000101",
-- "1010111100010110",
-- "1000110100010100",
-- "1100000000011101",
-- "0010100001000111",
-- "0111010100010011",
-- "0110101111010110",
-- "0001101010101111",
-- "1100100000111101",
-- "1011000101101111",
-- "1101010111000010",
-- "0000000111011100",
-- "0000100110000101",
-- "1111001111111111",
-- "1110111001010000",
-- "0001001111110100",
-- "0100100111100100",
-- "0101010100010101",
-- "0001011111010100",
-- "1011011110001111",
-- "1000000110100011",
-- "1010011000000011",
-- "0000100111000100",
-- "0101110111111101",
-- "0110010111010100",
-- "0010100101011011",
-- "1110011010010101",
-- "1101001010101001",
-- "1110101010000101",
-- "1111111111100011",
-- "1111000101011110",
-- "1101000100011100",
-- "1101000100001101",
-- "0000100100111000",
-- "0101010101001010",
-- "0111000001100010",
-- "0011011011111011",
-- "1100111000101010",
-- "1000011101000000",
-- "1001100001111011",
-- "1110110111100011",
-- "0011111001111010",
-- "0101000000000101",
-- "0010011110110100",
-- "1111101100011001",
-- "1111010011000000",
-- "0000101001101100",
-- "0000111010001100",
-- "1110100000111000",
-- "1011010100101000",
-- "1010111110100101",
-- "1111000100000001",
-- "0100111110100101",
-- "0111111001110011",
-- "0101001001111000",
-- "1110110001001001",
-- "1001110001001110",
-- "1001101110011010",
-- "1101110010100111",
-- "0001111100001010",
-- "0010111110111010",
-- "0001010110010000",
-- "0000000000111000",
-- "0000111100100000",
-- "0010110110010111",
-- "0010101000001110",
-- "1111000000000100",
-- "1010011011111000",
-- "1001001011011111",
-- "1101001000111100",
-- "0011101100001110",
-- "0111101110100101",
-- "0110001001111100",
-- "0000100101010010",
-- "1011101100011010",
-- "1010111100001011",
-- "1101101100111111",
-- "0000100000100000");--key8


-- "0110001001100001",
-- "0110110100100011",
-- "0010010010111110",
-- "1101110011011101",
-- "1101010101001100",
-- "1111011100001010",
-- "1111110111000101",
-- "1101010111101011",
-- "1011100100011110",
-- "1110010011000101",
-- "0100010010110110",
-- "0111110110000100",
-- "0101000000001101",
-- "1110001100100000",
-- "1001101110101100",
-- "1011000001101010",
-- "1111010110000111",
-- "0001100101110101",
-- "0000011001000000",
-- "1111001011001001",
-- "0001001100100000",
-- "0100110110011000",
-- "0101001111110100",
-- "0000010011010100",
-- "1001111011101011",
-- "1000001110011110",
-- "1100110011010001",
-- "0011000011000100",
-- "0101010010010001",
-- "0010110011001010",
-- "1111110110010010",
-- "0000000000000000",
-- "0001110101011011",
-- "0001001011110110",
-- "1100111111010011",
-- "1001010111000110",
-- "1011000011000011",
-- "0001100011110011",
-- "0111000110000001",
-- "0110101000110011",
-- "0001010001111110",
-- "1100101011010100",
-- "1100100101011101",
-- "1111000111101110",
-- "1111111000001100",
-- "1101110011111001",
-- "1100100011000010",
-- "1111100010011110",
-- "0101000100111100",
-- "0111100010010101",
-- "0011101011111010",
-- "1100101100010101",
-- "1000111100011011",
-- "1011001111101001",
-- "0000001011011000",
-- "0010011111100110",
-- "0001000111110111",
-- "1111101110010011",
-- "0001011010110001",
-- "0100011010111110",
-- "0100000100111001",
-- "1110111001101110",
-- "1001001100001000",
-- "1000101011011001",
-- "1110001001001110",
-- "0100011001100000",
-- "0101111011010100",
-- "0010101001101110",
-- "1111010001000111",
-- "1111010001011010",
-- "0001000000101011",
-- "0000010111111101",
-- "1100100110111010",
-- "1001110111110111",
-- "1100011001111001",
-- "0011000000111001",
-- "0111101101111100",
-- "0110000101010000",
-- "0000000001100011",
-- "1011100001111100",
-- "1100000001010010",
-- "1111000101111100",
-- "0000001100010101",
-- "1110011101001000",
-- "1101100011000110",
-- "0000100101011011",
-- "0101100000100100",
-- "0110111000010111",
-- "0010001101000111",
-- "1011010010111001",
-- "1000011110000100",
-- "1011110100010001",
-- "0001001111111000",
-- "0011011100001101",
-- "0001101101100110",
-- "0000000000000000",
-- "0001010100111010",
-- "0011110000010001",
-- "0010110110111111",
-- "1101101100101010",
-- "1000110011110111",
-- "1001011110111001",
-- "1111101001100010",
-- "0101101001100111",
-- "0110010001110111",
-- "0010001010111111",
-- "1110011100011001",
-- "1110011101110011",
-- "0000010010101101",
-- "1111110100111011",
-- "1100100100000100",
-- "1010101001110110",
-- "1101110100100010",
-- "0100010001001010",
-- "0111111110010100",
-- "0101001011100000",
-- "1110100110111101",
-- "1010011101110100",
-- "1011101101101000",
-- "1111011000010001",
-- "0000110000111111",
-- "1111001101111001",
-- "1110011110010101",
-- "0001010111011110",
-- "0101100101001100",
-- "0101111011111011",
-- "0000101010010001",
-- "1010000110011001",
-- "1000010110110001",
-- "1100101110010010",
-- "0010011110101100",
-- "0100010101010100",
-- "0010000101000010",
-- "1111111110010100",
-- "0000111101000010",
-- "0010111011101000",
-- "0001101100100110",
-- "1100110000111100",
-- "1000110011101111",
-- "1010100101011000",
-- "0001001101110100",
-- "0110101101001010",
-- "0110010010100100",
-- "0001010111110101",
-- "1101011100101001",
-- "1101101011011001",
-- "1111110000111100",
-- "1111100101001100",
-- "1100110101000101",
-- "1011100111110010",
-- "1111001100010011",
-- "0101001111100010",
-- "0111110110000010",
-- "0011111110111000",
-- "1101001000011001",
-- "1001100101001101",
-- "1011101110000110",
-- "1111111110010011",
-- "0001100010000010",
-- "0000000000000000",
-- "1111001111000000",
-- "0001110101110001",
-- "0101010100001010",
-- "0100110010001100",
-- "1111001010001010",
-- "1001001100000110",
-- "1000100111111000",
-- "1101111010100111",
-- "0011110001110111",
-- "0101000100101100",
-- "0010001010010010",
-- "1111101001001001",
-- "0000010110111001",
-- "0010000011001100",
-- "0000101011101111",
-- "1100001001110101",
-- "1001001010101100",
-- "1011111001110011",
-- "0010101111010011",
-- "0111011110110010",
-- "0101111011110101",
-- "0000010010111101",
-- "1100010111100010",
-- "1101000000011001",
-- "1111011111100111",
-- "1111101001010101",
-- "1101010110100010",
-- "1100101011100001",
-- "0000011010111100",
-- "0101111000011011",
-- "0111010101111100",
-- "0010100100010101",
-- "1011101100100100",
-- "1000111101100001",
-- "1100000100100100",
-- "0000110101101111",
-- "0010011010000101",
-- "0000101101001110",
-- "1111110000100000",
-- "0001111111010000",
-- "0100110000100111",
-- "0011100001010010",
-- "1101110011001110",
-- "1000100111110011",
-- "1001010000110001");--key9


-- "0101111010101100",
-- "0101101111000110",
-- "0001011001001111",
-- "1111100110100011",
-- "0010000101110101",
-- "0011011000010100",
-- "1111001011100111",
-- "1001010000001011",
-- "1000101011010001",
-- "1110001000011000",
-- "0010111101101101",
-- "0010011000000100",
-- "1111101011000000",
-- "0000110011110110",
-- "0101010000110111",
-- "0110011100111000",
-- "0001001110000100",
-- "1010110010000000",
-- "1001111010110010",
-- "1101111111001000",
-- "0000011000101000",
-- "1110001110111111",
-- "1100010101011100",
-- "1111110010110000",
-- "0110000000110110",
-- "0111101110011100",
-- "0010111010100100",
-- "1101100100111111",
-- "1101011001100001",
-- "0000001011110100",
-- "1111101110000100",
-- "1011010100001001",
-- "1001001100000110",
-- "1101100101111111",
-- "0100010111110100",
-- "0110010010001000",
-- "0010101001011000",
-- "1111101101110100",
-- "0001011010111011",
-- "0011110100011100",
-- "0001001011100000",
-- "1010110110110011",
-- "1000000011110110",
-- "1100000100101111",
-- "0001110000111001",
-- "0010101111111101",
-- "0000000001010101",
-- "1111110100100011",
-- "0100000001100101",
-- "0110111111011011",
-- "0011100001110101",
-- "1100100110100011",
-- "1001101010111111",
-- "1100101110110000",
-- "0000000110000111",
-- "1110111011001000",
-- "1100001001110001",
-- "1101111011010001",
-- "0100001010100011",
-- "0111111101011011",
-- "0100110111110011",
-- "1110111111110010",
-- "1101001100100000",
-- "1111101110100011",
-- "0000100011100011",
-- "1100101100011010",
-- "1001000000100010",
-- "1011011100011010",
-- "0010010100011111",
-- "0110001101010011",
-- "0011110110111101",
-- "0000001011011001",
-- "0000110000001000",
-- "0011110000100010",
-- "0010110111100010",
-- "1100111001010100",
-- "1000001101111000",
-- "1010010001101010",
-- "0000001010001011",
-- "0010110000010111",
-- "0000100011011101",
-- "1111001010001111",
-- "0010100011100101",
-- "0110110100011010",
-- "0101011101100101",
-- "1110110101010100",
-- "1010000101010000",
-- "1011100111000011",
-- "1111011110001010",
-- "1111100010001011",
-- "1100011011111000",
-- "1100011101010010",
-- "0001111111100101",
-- "0111011010100011",
-- "0110011101001101",
-- "0000101111111000",
-- "1101011001111111",
-- "1111001001111010",
-- "0001000001110110",
-- "1110001100110101",
-- "1001100001000110",
-- "1001110001101101",
-- "1111111110000001",
-- "0101011101100001",
-- "0100110101110000",
-- "0000111100100000",
-- "0000001111000010",
-- "0011010010000011",
-- "0100000101011011",
-- "1111001000110001",
-- "1001001000101100",
-- "1000111101001001",
-- "1110010011101101",
-- "0010010100001110",
-- "0001001000001000",
-- "1110111000001101",
-- "0001000011111110",
-- "0101111111111110",
-- "0110110100100011",
-- "0001001111011110",
-- "1011001010000000",
-- "1010110100000000",
-- "1110100101100110",
-- "1111111011011101",
-- "1101000100100000",
-- "1011100000111100",
-- "1111101111101010",
-- "0110001001011000",
-- "0111011110000101",
-- "0010101001011000",
-- "1110000101000010",
-- "1110100111101110",
-- "0001000111111000",
-- "1111101000100100",
-- "1010100111001010",
-- "1000110000100100",
-- "1101100100010110",
-- "0100000101000001",
-- "0101011010100000",
-- "0001111010011010",
-- "1111111111000000",
-- "0010100001110010",
-- "0100101111010111",
-- "0001010101001101",
-- "1010101101111101",
-- "1000010010001000",
-- "1100011010101101",
-- "0001011010100111",
-- "0001100101010110",
-- "1110111101011010",
-- "1111101110111001",
-- "0100101010111110",
-- "0111011110011100",
-- "0011100100011111",
-- "1100110100010111",
-- "1010011111101110",
-- "1101100100110010",
-- "0000000001001111",
-- "1101111001101110",
-- "1011001001100111",
-- "1101101010011110",
-- "0100010010110101",
-- "0111110001101000",
-- "0100011110001101",
-- "1111001100010000",
-- "1110010001110010",
-- "0000111000101110",
-- "0000110100100101",
-- "1100001000000000",
-- "1000011110101001",
-- "1011011000000010",
-- "0010001011010001",
-- "0101011100101000",
-- "0010111011011100",
-- "0000000011111100",
-- "0001101010011000",
-- "0100110100100000",
-- "0011001111101101",
-- "1100110010011111",
-- "1000010110111110",
-- "1010101101101100",
-- "0000000111010001",
-- "0001110001111111",
-- "1111010100110100",
-- "1110101101111010",
-- "0011000001101001",
-- "0111011000011000",
-- "0101100100010010",
-- "1110111010011111",
-- "1010110000111010",
-- "1100100110011000",
-- "1111110001101000",
-- "1110110000100111",
-- "1011010101101011",
-- "1011111101101110",
-- "0010000100000010",
-- "0111010100001100",
-- "0101111111111000",
-- "0000101001101100",
-- "1110010000001000",
-- "0000011011000111",
-- "0001101001000110",
-- "1101110110010110",
-- "1000111100000000",
-- "1001101000001110");--keyA


-- "0110000110111111",
-- "0101111011000001",
-- "0001010010010110",
-- "1110111111010100",
-- "0000111111001011",
-- "0010000101000000",
-- "1110001011011101",
-- "1001000100001000",
-- "1001100110101110",
-- "0000000101110110",
-- "0101011100010001",
-- "0100100011100111",
-- "0000101101100001",
-- "0000001001111010",
-- "0010111001101001",
-- "0010111111000011",
-- "1101101110011011",
-- "1000011110000000",
-- "1001101101100100",
-- "0000001010100111",
-- "0100011011010101",
-- "0010111011001010",
-- "0000001000100110",
-- "0001010110010000",
-- "0100101000101111",
-- "0011101011100110",
-- "1101011000111000",
-- "1000010101001000",
-- "1010001100101100",
-- "0000001101010101",
-- "0011000111111000",
-- "0001001000001101",
-- "1111100101111110",
-- "0010011111100101",
-- "0110000101101010",
-- "0100001000010111",
-- "1101001100110010",
-- "1000101010010001",
-- "1011000001110001",
-- "0000001101001111",
-- "0001100110110000",
-- "1111010001110110",
-- "1111000111101111",
-- "0011100001001011",
-- "0111001010101101",
-- "0100010100000111",
-- "1101001011100011",
-- "1001011100010100",
-- "1100001001001010",
-- "0000001001111000",
-- "1111111101110011",
-- "1101011111010110",
-- "1110101111100010",
-- "0100010110101011",
-- "0111110011101100",
-- "0100001110101110",
-- "1101010101111011",
-- "1010101000011000",
-- "1101011110001001",
-- "0000000011001000",
-- "1110010011011001",
-- "1011110111101011",
-- "1110011110011100",
-- "0100111100010110",
-- "0111111110001001",
-- "0011111001001000",
-- "1101101011111011",
-- "1100001001111011",
-- "1110111011010001",
-- "1111111001001111",
-- "1100101110000110",
-- "1010100001000100",
-- "1110010101000010",
-- "0101001111011000",
-- "0111101001011110",
-- "0011010101010000",
-- "1110001100110000",
-- "1101111011000101",
-- "0000011010101101",
-- "1111101100110111",
-- "1011010100010001",
-- "1001100000101001",
-- "1110010011001111",
-- "0101001110000100",
-- "0110110111000000",
-- "0010100101110110",
-- "1110110110110101",
-- "1111110100111111",
-- "0001110110100100",
-- "1111011110111101",
-- "1010001011101000",
-- "1000111010000111",
-- "1110011000100001",
-- "0100110111111100",
-- "0101101001111001",
-- "0001101110010010",
-- "1111100111111010",
-- "0001110000001100",
-- "0011001001010011",
-- "1111010000101111",
-- "1001011000111011",
-- "1000101111100100",
-- "1110100011110100",
-- "0100001101110110",
-- "0100000110111011",
-- "0000110010010010",
-- "0000011101001000",
-- "0011100101000110",
-- "0100001110000100",
-- "1111000011100110",
-- "1000111111100100",
-- "1001000001010110",
-- "1110110011101111",
-- "0011010001111011",
-- "0010010100001110",
-- "1111110101110000",
-- "0001010011001110",
-- "0101001100100001",
-- "0101000000111101",
-- "1110111000111100",
-- "1001000001011110",
-- "1001101110000101",
-- "1111000110101100",
-- "0010000111011101",
-- "0000011000110110",
-- "1110111100011101",
-- "0010000110101100",
-- "0110100000000010",
-- "0101011111010000",
-- "1110110010000111",
-- "1001011110110110",
-- "1010110010101100",
-- "1111011010111101",
-- "0000110010110001",
-- "1110011100011010",
-- "1110001001110010",
-- "0010110100000110",
-- "0111011010011100",
-- "0101100111100100",
-- "1110110000010000",
-- "1010010110001110",
-- "1100001010101111",
-- "1111101110111010",
-- "1111011000111011",
-- "1100100110011111",
-- "1101100000100110",
-- "0011011000001011",
-- "0111111000000010",
-- "0101011001111001",
-- "1110110100001100",
-- "1011100100011111",
-- "1101110000100111",
-- "0000000001000011",
-- "1101111111011010",
-- "1010111110010011",
-- "1101000011000001",
-- "0011110000001100",
-- "0111110110111010",
-- "0100110111100111",
-- "1110111110010101",
-- "1101000101000101",
-- "1111011101111001",
-- "0000010000001101",
-- "1100101011110101",
-- "1001101010001011",
-- "1100110010010101",
-- "0011111010000100",
-- "0111010111000011",
-- "0100000011010011",
-- "1111001110100101",
-- "1110110010001110",
-- "0001001011110110",
-- "0000011011100010",
-- "1011100011100011",
-- "1000101111001000",
-- "1100101110111110",
-- "0011110100100100",
-- "0110011010010100",
-- "0011000000100110",
-- "1111100100011000",
-- "0000100101010100",
-- "0010110011101110",
-- "0000100010101000",
-- "1010101011010011",
-- "1000010000101100",
-- "1100111000011111",
-- "0011011111011000",
-- "0101000100010110",
-- "0001110011111101",
-- "1111111110101010",
-- "0010010111010100",
-- "0100001111010010",
-- "0000100101011110",
-- "1010000110111101",
-- "1000010000100101",
-- "1101001101101001",
-- "0010111011010001",
-- "0011011010011000",
-- "0000100010010101",
-- "0000011011111010",
-- "0100000001001100",
-- "0101011001000101",
-- "0000100100011100",
-- "1001111001001100",
-- "1000101110100111");--keyB

-- "0110010100010000",
-- "0110000100101010",
-- "0001000001111000",
-- "1110001000110100",
-- "1111101101001011",
-- "0000111000100100",
-- "1101101110101111",
-- "1001110100111010",
-- "1011100011011010",
-- "0010100111010010",
-- "0111100001011000",
-- "0101001011111011",
-- "1111010111011011",
-- "1101000110111100",
-- "1111001101110110",
-- "0000001001010101",
-- "1101000010000011",
-- "1010011100111011",
-- "1101110100100001",
-- "0100111001011101",
-- "0111111000010101",
-- "0011100100011001",
-- "1101011111000101",
-- "1100010000000000",
-- "1111000000001111",
-- "1111110001011100",
-- "1100111001010001",
-- "1011101001000110",
-- "0000001011010001",
-- "0110100100011101",
-- "0111010100101011",
-- "0001011000110000",
-- "1011101001101100",
-- "1011110001101110",
-- "1111001100001110",
-- "1111110011010111",
-- "1101001111011001",
-- "1101001010101111",
-- "0010010100000100",
-- "0111011011110110",
-- "0101111010000000",
-- "1110111001100001",
-- "1010001001001010",
-- "1011110110101111",
-- "1111110100011011",
-- "0000001011101110",
-- "1101111010011101",
-- "1110110001001101",
-- "0011111110011011",
-- "0111011010011111",
-- "0011110011011110",
-- "1100011010110001",
-- "1001001101101001",
-- "1100100100011110",
-- "0000110101100001",
-- "0000110010001000",
-- "1110101101100100",
-- "0000001100110000",
-- "0100111111010001",
-- "0110100011001010",
-- "0001010010010000",
-- "1010010001001111",
-- "1001000010110111",
-- "1101111001111001",
-- "0010000110100011",
-- "0001011010110011",
-- "1111011011011110",
-- "0001010001000001",
-- "0101010010010100",
-- "0100111111111000",
-- "1110101010111111",
-- "1000101111010011",
-- "1001101110000001",
-- "1111101111001010",
-- "0011011010010100",
-- "0001111000111000",
-- "1111111001000000",
-- "0001110110111010",
-- "0100111010011001",
-- "0011000000010000",
-- "1100010010110100",
-- "1000000010001010",
-- "1011001100110000",
-- "0001110110100011",
-- "0100100001011100",
-- "0010000000111100",
-- "1111111111001100",
-- "0001111101011011",
-- "0100000000100011",
-- "0000110110111011",
-- "1010011100010110",
-- "1000001111111100",
-- "1101010101001010",
-- "0011111110010110",
-- "0101001101001001",
-- "0001101011011000",
-- "1111101100100010",
-- "0001101001100011",
-- "0010110010001100",
-- "1110110110101010",
-- "1001010100111110",
-- "1001010110101111",
-- "1111110111000110",
-- "0101110011011011",
-- "0101010001110000",
-- "0000110101111101",
-- "1111000101010100",
-- "0001000100111111",
-- "0001011110101100",
-- "1101001111100001",
-- "1001000011000111",
-- "1011001100111010",
-- "0010011110011001",
-- "0111000100001101",
-- "0100101001000001",
-- "1111100100101010",
-- "1110010010110000",
-- "0000011100000111",
-- "0000010100100111",
-- "1100001100100101",
-- "1001100101011111",
-- "1101100010100010",
-- "0100110101101111",
-- "0111100011011010",
-- "0011010011011011",
-- "1110000001010110",
-- "1101100001010101",
-- "1111111011100110",
-- "1111011111010101",
-- "1011110010011110",
-- "1010110011101010",
-- "0000000011110001",
-- "0110101001101111",
-- "0111001010010000",
-- "0001011000100111",
-- "1100011010010011",
-- "1100111110100000",
-- "1111101101110100",
-- "1111000101001100",
-- "1011111111000010",
-- "1100011111100010",
-- "0010011011110110",
-- "0111101011110101",
-- "0101111001101101",
-- "1111000110011110",
-- "1011000000000110",
-- "1100110110000100",
-- "1111111000111001",
-- "1111000110100101",
-- "1100101010001100",
-- "1110010111110100",
-- "0100011000000011",
-- "0111110100010001",
-- "0011111010011110",
-- "1100101111010101",
-- "1010000010110101",
-- "1101001111110110",
-- "0000011101010111",
-- "1111011110001100",
-- "1101100111100001",
-- "0000001010110011",
-- "0101101010011010",
-- "0111000011001111",
-- "0001011011111100",
-- "1010100111010100",
-- "1001101111011101",
-- "1110001101111111",
-- "0001010110000010",
-- "0000000010001110",
-- "1110101000110100",
-- "0001101001001010",
-- "0110001011100011",
-- "0101100000110000",
-- "1110110001111101",
-- "1001000001010101",
-- "1010001101011001",
-- "1111101100001000",
-- "0010011000101001",
-- "0000100110010101",
-- "1111100000101000",
-- "0010101000001101",
-- "0101111011100001",
-- "0011011011010010",
-- "1100010010000010",
-- "1000001100001100",
-- "1011011101000101",
-- "0001011111110001",
-- "0011010111101110",
-- "0000111110001010",
-- "0000000100100110",
-- "0011000011010111",
-- "0101000001010110",
-- "0001000101100001",
-- "1010010000001101",
-- "1000010000010110",
-- "1101010111100001",
-- "0011011001101100",
-- "0100000100111101",
-- "0000111111110001",
-- "0000001111011000",
-- "0010111100011111",
-- "0011101001101101",
-- "1110110011100000",
-- "1000111100001000",
-- "1001001110011110");--keyC

-- "0111111111111111",
-- "0111111111111111",
-- "0001001100100000",
-- "1010001010011010",
-- "1100110100111100",
-- "0000001101001111",
-- "1100010010101110",
-- "1000000000000000",
-- "1100000011001011",
-- "0111111111111111",
-- "0111111111111111",
-- "0110101110000000",
-- "1000000000000000",
-- "1000000000000000",
-- "1011000100001010",
-- "0010100011101001",
-- "0001011110010110",
-- "1110010000111001",
-- "0010011011011010",
-- "0111111111111111",
-- "0111111111111111",
-- "1100010001100010",
-- "1000000000000000",
-- "1000000000000000",
-- "0001111010011010",
-- "0111111111111111",
-- "0110100100111010",
-- "1111111000111111",
-- "0000010111100100",
-- "0100001011001101",
-- "0000101100101011",
-- "1000000000000000",
-- "1000000000000000",
-- "1101000001110111",
-- "0111111111111111",
-- "0111111111111111",
-- "0011110011111100",
-- "1001100001001100",
-- "1001111000001110",
-- "1111001101000010",
-- "1110101011100011",
-- "1001100000110111",
-- "1010111101101010",
-- "0110001101100011",
-- "0111111111111111",
-- "0111111111111111",
-- "1010001000011011",
-- "1000000000000000",
-- "1000001000101101",
-- "0010010001001111",
-- "0100001101101101",
-- "0000000100110100",
-- "0000101100010100",
-- "0111100011110100",
-- "0111111111111111",
-- "1111001100111100",
-- "1000000000000000",
-- "1000000000000000",
-- "1111001100111110",
-- "0111111111111111",
-- "0111111111111111",
-- "0001000100110101",
-- "1110000110100100",
-- "0001101110110001",
-- "0001100110111001",
-- "1001011010100110",
-- "1000000000000000",
-- "1010011101110111",
-- "0111111111111111",
-- "0111111111111111",
-- "0110110010100001",
-- "1001111111001110",
-- "1000000000000000",
-- "1101001111011101",
-- "0000010000000111",
-- "1100010110101001",
-- "1010111110011010",
-- "0011010110001000",
-- "0111111111111111",
-- "0111111111111111",
-- "1100111010101001",
-- "1000000000000000",
-- "1000000000000000",
-- "0000111010001100",
-- "0110010111000000",
-- "0010100111101110",
-- "1111111110000000",
-- "0100100110010111",
-- "0111111111111111",
-- "0001101010011001",
-- "1000000000000000",
-- "1000000000000000",
-- "1100001100010101",
-- "0111111111111111",
-- "0111111111111111",
-- "0011001011110101",
-- "1100101100100011",
-- "1110110110011100",
-- "0001011010010010",
-- "1100001101000110",
-- "1000000000000000",
-- "1000101010100001",
-- "0110100011001100",
-- "0111111111111111",
-- "0111111111111111",
-- "1011100000101010",
-- "1000000000000000",
-- "1010100110000101",
-- "0000110010010010",
-- "1111010010011111",
-- "1100000101000000",
-- "0001000000010111",
-- "0111111111111111",
-- "0111111111111111",
-- "1111111100000010",
-- "1000000000000000",
-- "1000000000000000",
-- "1110101010011001",
-- "0111100110110001",
-- "0101100010101011",
-- "0000010110111001",
-- "0001111001010100",
-- "0110100110011101",
-- "0011010100001111",
-- "1000000000000000",
-- "1000000000000000",
-- "1001010011000000",
-- "0111111111111111",
-- "0111111111111111",
-- "0101111011010010",
-- "1100010110010101",
-- "1011111100001101",
-- "0000001000110001",
-- "1110011010010110",
-- "1000000000000000",
-- "1000000000000000",
-- "0011100010011001",
-- "0111111111111111",
-- "0111111111111111",
-- "1101111000010000",
-- "1000000000000000",
-- "1000000000000000",
-- "0000001101001001",
-- "0001111001111001",
-- "1110000111010010",
-- "1111100000111101",
-- "0111111111111111",
-- "0111111111111111",
-- "0010110010000000",
-- "1000000000000000",
-- "1000000000000000",
-- "1011110101100111",
-- "0111110001100011",
-- "0111111111111111",
-- "0001110011011110",
-- "1111110101000000",
-- "0011111111111100",
-- "0011111100000010",
-- "1010100010111001",
-- "1000000000000000",
-- "1000000000000000",
-- "0110000011000101",
-- "0111111111111111",
-- "0111111111111111",
-- "1101000111010011",
-- "1001011010010101",
-- "1101111101111101",
-- "1111101110101010",
-- "1010100111100011",
-- "1000001011110001",
-- "0000110001000101",
-- "0111111111111111",
-- "0111111111111111",
-- "0000110001001101",
-- "1000000000000000",
-- "1000000000000000",
-- "1110100101101110",
-- "0011110101010000",
-- "0000110010110011",
-- "1111000101000100",
-- "0101000111010100",
-- "0111111111111111",
-- "0101000011100001",
-- "1000000000000000",
-- "1000000000000000",
-- "1000110100110100",
-- "0110110101100001",
-- "0111111111111111",
-- "0100000110110011",
-- "1110101100000010",
-- "0001000100011010",
-- "0011011100100001",
-- "1101001110011010",
-- "1000000000000000",
-- "1000000000000000",
-- "0011000111010000",
-- "0111111111111111",
-- "0111111111111111",
-- "1110111000111010",
-- "1000000000000000",
-- "1011001101010110",
-- "1111111110001111",
-- "1101100000110111",
-- "1001100011111110",
-- "1110100111101110");--keyD

begin
process(clk_5mhz,rst,en)
begin
		
	if(clk_5mhz'event and clk_5mhz = '1')  then 			
		if rst = '1' then 			
			ram_out <=(others=>'0');			
		elsif en='1' then
			ram_out <= ram1(conv_integer(addr));
		else--changed
			ram_out <=(others=>'0');		
	end if;
end if;	
end process;
end Behavioral;

