----------------------------------------------------------------------------------
-- Company: CEM Solutions
-- Engineer: viru jawoor
-- 
-- Create Date:    17:30:26 05/20/2008 
-- Design Name:    RINGING TONE 
-- Module Name:    RAM- Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: SINE WAVE At 770Hz
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity SIG_RAM is
    Port ( clk_5mhz : in  STD_LOGIC;
           rst : in  STD_LOGIC;
           en : in  STD_LOGIC;
		   addr : in std_logic_vector(7 downto 0);
           ram_out : out  STD_LOGIC_vector(15 downto 0));
end SIG_RAM;

architecture Behavioral of SIG_RAM is

type ram is array  (0 to 204)of std_logic_vector (15 downto 0);
constant ram1 : ram :=(--"0001001000110010",
--"0001110111101111",
--"0001111100001110",
--"0001010100101001",
--"0000001111000011",
--"1111000100000111",
--"1110001110011010",
--"1110000001000001",
--"1110100000101010",
--"1111100010001000",
--"0000101110001100",
--"0001101001110111",
--"0010000000000000",
--"0001101000101110",
--"0000101100010011",
--"1111100000001011",
--"1110011111010101",
--"1110000000110001",
--"1110001111010111",
--"1111000101111001",
--"0000010001000011",
--"0001010110001001",
--"0001111100101100",
--"0001110111000001",
--"0001000111000111",
--"1111111101111111",
--"1110110101100101",
--"1110000111100100",
--"1110000100010010",
--"1110101100111000",
--"1111110010111101",
--"0000111101101011",
--"0001110010100000",
--"0001111110101110",
--"0001011110000000",
--"0000011011111011",
--"1111001111111101",
--"1110010101000001",
--"1110000000000010",
--"1110011000011101",
--"1111010101100110",
--"0000100001110010",
--"0001100001111111",
--"0001111111011100",
--"0001101111101011",
--"0000111000010100",
--"1111101100111110",
--"1110101000011000",
--"1110000010111000",
--"1110001001110000",
--"1110111010100100",
--"0000000100000001",
--"0001001100000011",
--"0001111001000110",
--"0001111011001100",
--"0001010001100110",
--"0000001011000011",
--"1111000000100101",
--"1110001100100111",
--"1110000001100101",
--"1110100011011001",
--"1111100110000011",
--"0000110001111010",
--"0001101100000101",
--"0001111111111010",
--"0001100110010111",
--"0000101000100001",
--"1111011100010011",
--"1110011100101111",
--"1110000000011001",
--"1110010001010100",
--"1111001001100000",
--"0000010101000001",
--"0001011001000101",
--"0001111101100011",
--"0001110101011110",
--"0001000011101111",
--"1111111001111110",
--"1110110010010110",
--"1110000110010001",
--"1110000101010111",
--"1110101111111110",
--"1111110110111101",
--"0001000001001010",
--"0001110100010000",
--"0001111110000110",
--"0001011011001110",
--"0000010111111111",
--"1111001100010000",
--"1110010010110111",
--"1110000000001100",
--"1110011010110111",
--"1111011001011010",
--"0000100101101001",
--"0001100100100001",
--"0001111111110000",
--"0001101101101010",
--"0000110100101011",
--"1111101001000000",
--"1110100101011111",
--"1110000010000101",
--"1110001011010110",
--"1110111101111111",
--"0000001000000010",
--"0001001111010000",
--"0001111010010110",
--"0001111010000011",
--"0001001110011101",
--"0000000111000010",
--"1110111101001000",
--"1110001010111100",
--"1110000010010001",
--"1110100110001101",
--"1111101010000000",
--"0000110101100110",
--"0001101110001011",
--"0001111111101100",
--"0001100011111001",
--"0000100100101011",
--"1111011000011101",
--"1110011010010000",
--"1110000000001001",
--"1110010011011001",
--"1111001101001011",
--"0000011000111110",
--"0001011011111011",
--"0001111110010001",
--"0001110011110100",
--"0001000000010011",
--"1111110101111101",
--"1110101111001100",
--"1110000101000101",
--"1110000110100101",
--"1110110011001001",
--"1111111010111110",
--"0001000100100101",
--"0001110101111000",
--"0001111101010110",
--"0001011000010111",
--"0000010100000010",
--"1111001000100110",
--"1110010000110100",
--"1110000000011111",
--"1110011101011000",
--"1111011101010000",
--"0000101001011110",
--"0001100110111101",
--"0001111111111100",
--"0001101011100010",
--"0000110000111111",
--"1111100101000100",
--"1110100010101100",
--"1110000001011011",
--"1110001101000011",
--"1111000001011101",
--"0000001100000011",
--"0001010010010111",
--"0001111011011110",
--"0001111000110001",
--"0001001011001111",
--"0000000011000001",
--"1110111001101110",
--"1110001001010111",
--"1110000011000101",
--"1110101001000111",
--"1111101101111110",
--"0000111001001110",
--"0001110000001011",
--"0001111111010101",
--"0001100001010101",
--"0000100000110100",
--"1111010100101001",
--"1110010111110111",
--"1110000000000001",
--"1110010101100101",
--"1111010000111000",
--"0000011100111010",
--"0001011110101011",
--"0001111110110111",
--"0001110010000011",
--"0000111100110010",
--"1111110001111101",
--"1110101100000111",
--"1110000100000001",
--"1110000111111010",
--"1110110110011010",
--"1111111111000000",
--"0001000111111101",
--"0001110111011000",
--"0001111100011110",
--"0001010101011010",
--"0000010000000011",
--"1111000101000000",
--"1110001110111000",
--"1110000000111001",
--"1110011111111111",
--"1111100001001001",
--"0000101101010000",
--"0001101001010011",
--"0010000000000000",
--"0001101001010011",
--"0000101101010000",
--"1111100001001001",
--"1110011111111111",
--"1110000000111001");

"0011101010101101",
"0010111011011100",
"1110101010111111",
"1100000000101011",
"1110001001000110",
"0010100000011000",
"0011110110111111",
"0000100100110111",
"1100100110011110",
"1100101101011010",
"0000110001010110",
"0011111010000001",
"0010010110010100",
"1101111110000010",
"1100000001111001",
"1110110111000010",
"0011000011110101",
"0011100101010111",
"1111110011010110",
"1100010000100010",
"1101001101011010",
"0001100000110110",
"0011111111111100",
"0001101011100011",
"1101010101111101",
"1100001100101010",
"1111100111101101",
"0011011111111101",
"0011001011001001",
"1111000010010010",
"1100000011100101",
"1101110100001000",
"0010001100101110",
"0011111100010000",
"0000111100101111",
"1100110100010000",
"1100100000100011",
"0000011001010011",
"0011110011101010",
"0010101001010011",
"1110010011100011",
"1100000000000110",
"1110100000000101",
"0010110011010100",
"0011101111000111",
"0000001011101010",
"1100011010001100",
"1100111100110100",
"0001001001111011",
"0011111110001110",
"0010000001000110",
"1101101000111000",
"1100000110001101",
"1111001111101001",
"0011010011001011",
"0011011001000000",
"1111011010001001",
"1100001000110000",
"1101100000011010",
"0001110111110011",
"0011111111010000",
"0001010100000100",
"1101000011111000",
"1100010101101101",
"0000000001000000",
"0011101011000111",
"0010111010110000",
"1110101010000011",
"1100000000100110",
"1110001001111111",
"0010100001001010",
"0011110110101110",
"0000100011111000",
"1100100101111100",
"1100101101111111",
"0000110010010110",
"0011111010001110",
"0010010101100000",
"1101111101001011",
"1100000010000001",
"1110111000000000",
"0011000100011111",
"0011100100111010",
"1111110010010101",
"1100010000001011",
"1101001110001001",
"0001100001110010",
"0011111111111101",
"0001101010101000",
"1101010101001101",
"1100001100111110",
"1111101000101101",
"0011100000011100",
"0011001010100010",
"1111000001010100",
"1100000011011010",
"1101110100111110",
"0010001101100100",
"0011111100000101",
"0000111011110001",
"1100110011101001",
"1100100001000010",
"0000011010010011",
"0011110011111110",
"0010101000100011",
"1110010010101001",
"1100000000001000",
"1110100001000001",
"0010110100000001",
"0011101110110000",
"0000001010101010",
"1100011001110000",
"1100111101011110",
"0001001010111001",
"0011111110010110",
"0010000000001111",
"1101101000000100",
"1100000110011100",
"1111010000101000",
"0011010011101111",
"0011011000011110",
"1111011001001001",
"1100001000100000",
"1101100001001101",
"0001111000101011",
"0011111111001011",
"0001010011000111",
"1101000011001101",
"1100010110000111",
"0000000010000001",
"0011101011100000",
"0010111010000100",
"1110101001000110",
"1100000000100010",
"1110001010111001",
"0010100001111100",
"0011110110011100",
"0000100010111000",
"1100100101011010",
"1100101110100011",
"0000110011010101",
"0011111010011100",
"0010010100101011",
"1101111100010011",
"1100000010001001",
"1110111000111110",
"0011000101001000",
"0011100100011110",
"1111110001010101",
"1100001111110101",
"1101001110110111",
"0001100010101101",
"0011111111111110",
"0001101001101110",
"1101010100011101",
"1100001101010010",
"1111101001101101",
"0011100000111010",
"0011001001111010",
"1111000000010101",
"1100000011010000",
"1101110101110100",
"0010001110011001",
"0011111011111010",
"0000111010110010",
"1100110011000011",
"1100100001100010",
"0000011011010011",
"0011110100010001",
"0010100111110010",
"1110010001101111",
"1100000000001010",
"1110100001111101",
"0010110100101111",
"0011101110011001",
"0000001001101010",
"1100011001010100",
"1100111110001000",
"0001001011110110",
"0011111110011101",
"0001111111010111",
"1101100111010001",
"1100000110101010",
"1111010001100111",
"0011010100010011",
"0011010111111100",
"1111011000001010",
"1100001000010000",
"1101100001111111",
"0001111001100100",
"0011111111000110",
"0001010010001010",
"1101000010100001",
"1100010110100001",
"0000000011000001",
"0011101011111001",
"0010111001011000",
"1110101000001010",
"1100000000011110",
"1110001011110010",
"0010100010101110",
"0011110110001011",
"0000100001111000",
"1100100100111001",
"1100101111001001");




begin
process(clk_5mhz,rst,en)
begin
		
	if(clk_5mhz'event and clk_5mhz = '0')  then 			
		if rst = '1' then 			
			ram_out <=(others=>'0');			
		elsif en='1' then
			ram_out <= ram1(conv_integer(addr));
		else--changed
		ram_out <=(others=>'0');		
	end if;
end if;	
end process;
end Behavioral;

